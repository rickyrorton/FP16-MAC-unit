module control (data_in,store_num,mac_clk,result);
    
endmodule