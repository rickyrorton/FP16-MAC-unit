//-----------------------------------------------------------
// File: fpu_tb.v
// FPU Test Bench
//-----------------------------------------------------------
`timescale 1 ns/100 ps
module fpu_tb ();
 //----------------------------------------------------------
 // inputs to the DUT are reg type
 reg clock;
 reg [31:0] a, b;
 reg [1:0] op;
 reg [31:0] correct;
 //----------------------------------------------------------
 // outputs from the DUT are wire type
 wire [31:0] out;
 wire [49:0] pro;
 //----------------------------------------------------------
 // instantiate the Device Under Test (DUT)
 // using named instantiation
 fpu U1 (
          .clk(clock),
          .A(a),
          .B(b),
          .opcode(op),
          .O(out)
        );
 //----------------------------------------------------------
 // create a 10Mhz clock
 always
 #100 clock = ~clock; // every 100 nanoseconds invert
 //----------------------------------------------------------
 // initial blocks are sequential and start at time 0
 initial
 begin
 $dumpfile("fpu_tb.vcd");
 $dumpvars(0,clock, a, b, op, out);
 clock = 0;a = 16'b00111110001010001100000000000000;
b = 16'b00111010000001011000000000000000;
a = 16'b01000101011111011100000000000000;
b = 16'b11000101010101000110000000000000;
a = 16'b01000111010001111110000000000000;
b = 16'b10110111101111001000000000000000;
a = 16'b11000001000110001110000000000000;
b = 16'b11000000110001001010000000000000;
a = 16'b11000000010101110000000000000000;
b = 16'b11000000001010111100000000000000;
a = 16'b10111011010011001100000000000000;
b = 16'b00111010011010011100000000000000;
a = 16'b10111101100101011010000000000000;
b = 16'b01000000001000100000000000000000;
a = 16'b10111010100011101000000000000000;
b = 16'b10111001111101000110000000000000;
a = 16'b00111011101011100110000000000000;
b = 16'b00111101110000100000000000000000;
a = 16'b11000100100010001100000000000000;
b = 16'b01000101000010001000000000000000;
$display ("Done.");
$finish;
 // stop the simulation
 end

endmodule